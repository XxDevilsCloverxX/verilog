module Hello;
// This is a comment
initial begin
$display("Hello World");
$finish;
end
endmodule